library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ramp_gen is
	generic(
	  COUNT_NBITS: integer := 18;     -- number of bits of the counter
  	COUNT_MOD: integer := 200000;		-- mod-n
		DATA_BITS: integer := 12);			-- number of bits for the data
  port(
    aclk       			: in    std_logic;
		aresetn					: in 		std_logic;
		data_i					: in 		std_logic_vector(DATA_BITS-1 downto 0);
		data_o				: out 	std_logic_vector(DATA_BITS-1 downto 0);
		pwm_o				: out		std_logic;
		led_o		: out 	std_logic);
end ramp_gen;

architecture rtl of ramp_gen is
  signal cnt_reg, cnt_next	: unsigned(COUNT_NBITS-1 downto 0);
  signal in_reg, in_next	: unsigned(DATA_BITS-1 downto 0);
  signal r_reg, r_next	: unsigned(DATA_BITS-1 downto 0);
  signal out_reg, out_next	: unsigned(DATA_BITS-1 downto 0);
	signal buff_reg, buff_next			: std_logic;
	signal max_tick			: std_logic;

begin
	-- Drive inputs
	in_next	<= unsigned(data_i);

	--registers
 	process (aclk)
 	begin
    if rising_edge(aclk) then
      if (aresetn = '0') then
    	  cnt_reg 	<= (others => '0');
    	  in_reg 		<= (others => '0');
    	  out_reg 	<= (others => '0');
    	  r_reg		 	<= (others => '0');
    	  buff_reg 	<= '0';
      else
     	  cnt_reg 	<= cnt_next;
     	  r_reg 		<= r_next;
     	  buff_reg 		<= buff_next;
     	  in_reg 		<= in_next;
     	  out_reg 	<= out_next;
      end if;
    end if;
 	end process;
	--next-state logic for counter
	cnt_next	<= 	(others => '0') when cnt_reg = (COUNT_MOD-1) else
          				cnt_reg + 1;

	buff_next <= '1' when (r_reg < out_reg) else '0';          		

	r_next <= r_reg + 1;          		

	--output logic
	max_tick <= '1' when cnt_reg = (COUNT_MOD-1) else '0';

	process(max_tick, in_reg, out_reg)
	begin
		if (max_tick = '1') then
			if (in_reg > out_reg) then			
				out_next <= out_reg + 1;
			elsif (in_reg < out_reg) then
				out_next <= out_reg - 1;
			else
				out_next <= out_reg;	-- default
			end if;
		else
			out_next <= out_reg;
		end if;
	end process;
	
	--next-state logic for output
	data_o	<= std_logic_vector(out_reg);
	led_o <= 	'0' when (out_reg = 0) else
						'1';
	pwm_o <= buff_reg;

end rtl;
